`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/06/2018 03:17:58 PM
// Design Name: 
// Module Name: sub4hex
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

//declare inputs and outputs
module sub4hex(
  input [3:0] A,
  input [3:0] B,
  output [3:0] Sum,
  output [6:0] segs7,
  output [3:0] anodes
  );

  wire of_s,c_msb;
  wire negB;
  
 
endmodule
